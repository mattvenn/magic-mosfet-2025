MOSFET Simulation
* this file edited to remove everything not in tt lib
.lib "/foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.include mosfet.spice

* instantiate the extracted MOSFET
Xmosfet GATE DRAIN VGND mosfet

* set gnd and power
Vgnd VGND 0 0
Vdd VPWR VGND 1.8
Vsubs VSUBS 0 0

* create a resistor between the MOSFET drain and VPWR
R VPWR DRAIN 10k

* create pulse
Vin GATE VGND pulse(0 1.8 1p 10p 10p 1n 2n)
.tran 10p 2n 0

.control
run
set color0 = white
set color1 = black
plot GAIN DRAIN
.endc

.end
