magic
tech sky130A
timestamp 1752846654
<< nmos >>
rect 40 0 55 65
<< ndiff >>
rect 0 0 40 65
rect 55 0 95 65
<< poly >>
rect 40 65 55 105
rect 40 -45 55 0
<< labels >>
flabel poly 40 65 55 105 0 FreeSans 80 0 0 0 gate
port 1 nsew
flabel ndiff 0 0 40 65 0 FreeSans 80 0 0 0 drain
port 2 nsew
flabel ndiff 55 0 95 65 0 FreeSans 80 0 0 0 source
port 3 nsew
<< end >>
